	component unsaved is
		port (
			clk_50_clk    : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component unsaved;

	u0 : component unsaved
		port map (
			clk_50_clk    => CONNECTED_TO_clk_50_clk,    -- clk_50.clk
			reset_reset_n => CONNECTED_TO_reset_reset_n  --  reset.reset_n
		);

