
module unsaved (
	clk_50_clk,
	reset_reset_n);	

	input		clk_50_clk;
	input		reset_reset_n;
endmodule
